VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BATCHARGERctr
  CLASS BLOCK ;
  ORIGIN -19.5 -7.1 ;
  FOREIGN BATCHARGERctr 19.5 7.1 ;
  SIZE 83.8 BY 41.8 ;
  SYMMETRY X Y R90 ;
  PIN dvdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME3 ;
        RECT 19.5 45.9 19.7 46.1 ;
    END
  END dvdd
  PIN dgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME3 ;
        RECT 19.5 45.1 19.7 45.3 ;
    END
  END dgnd
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME2 ;
        RECT 21.1 7.1 21.3 7.3 ;
    END
  END clk
  PIN iend
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 19.5 19.9 19.7 20.1 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 19.5 19.7 19.7 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 19.1 19.7 19.3 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 18.7 19.7 18.9 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 18.3 19.7 18.5 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 17.9 19.7 18.1 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 17.5 19.7 17.7 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 17.1 19.7 17.3 ;
    END
  END iend
  PIN vcutoff
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 19.5 39.9 19.7 40.1 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 39.5 19.7 39.7 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 39.1 19.7 39.3 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 38.7 19.7 38.9 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 38.3 19.7 38.5 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 37.9 19.7 38.1 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 37.5 19.7 37.7 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 37.1 19.7 37.3 ;
    END
  END vcutoff
  PIN vpreset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 19.5 35.9 19.7 36.1 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 35.5 19.7 35.7 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 35.1 19.7 35.3 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 34.7 19.7 34.9 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 34.3 19.7 34.5 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 33.9 19.7 34.1 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 33.5 19.7 33.7 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 33.1 19.7 33.3 ;
    END
  END vpreset
  PIN tmax
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 19.5 23.9 19.7 24.1 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 23.5 19.7 23.7 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 23.1 19.7 23.3 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 22.7 19.7 22.9 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 22.3 19.7 22.5 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 21.9 19.7 22.1 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 21.5 19.7 21.7 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 21.1 19.7 21.3 ;
    END
  END tmax
  PIN tempmax
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 19.5 27.9 19.7 28.1 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 27.5 19.7 27.7 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 27.1 19.7 27.3 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 26.7 19.7 26.9 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 26.3 19.7 26.5 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 25.9 19.7 26.1 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 25.5 19.7 25.7 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 25.1 19.7 25.3 ;
    END
  END tempmax
  PIN tempmin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 19.5 31.9 19.7 32.1 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 31.5 19.7 31.7 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 31.1 19.7 31.3 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 30.7 19.7 30.9 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 30.3 19.7 30.5 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 29.9 19.7 30.1 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 29.5 19.7 29.7 ;
    END
    PORT
      LAYER ME3 ;
        RECT 19.5 29.1 19.7 29.3 ;
    END
  END tempmin
  PIN vbat
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 39.9 7.1 40.1 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 40.3 7.1 40.5 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 40.7 7.1 40.9 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 41.1 7.1 41.3 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 41.5 7.1 41.7 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 41.9 7.1 42.1 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 42.3 7.1 42.5 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 42.7 7.1 42.9 7.3 ;
    END
  END vbat
  PIN vmonem
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 51.9 7.1 52.1 7.3 ;
    END
  END vmonem
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 23.5 7.1 23.7 7.3 ;
    END
  END en
  PIN rstz
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 21.9 7.1 22.1 7.3 ;
    END
  END rstz
  PIN vtok[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 19.5 15.9 19.7 16.1 ;
    END
  END vtok[0]
  PIN ibat
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 43.9 7.1 44.1 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 44.3 7.1 44.5 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 44.7 7.1 44.9 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 45.1 7.1 45.3 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 45.5 7.1 45.7 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 45.9 7.1 46.1 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 46.3 7.1 46.5 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 46.7 7.1 46.9 7.3 ;
    END
  END ibat
  PIN tbat
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 47.9 7.1 48.1 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 48.3 7.1 48.5 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 48.7 7.1 48.9 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 49.1 7.1 49.3 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 49.5 7.1 49.7 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 49.9 7.1 50.1 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 50.3 7.1 50.5 7.3 ;
    END
    PORT
      LAYER ME2 ;
        RECT 50.7 7.1 50.9 7.3 ;
    END
  END tbat
  PIN cc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 103.1 11.9 103.3 12.1 ;
    END
  END cc
  PIN tc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 103.1 10.3 103.3 10.5 ;
    END
  END tc
  PIN cv
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 103.1 11.1 103.3 11.3 ;
    END
  END cv
  PIN imonem
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 53.1 7.1 53.3 7.3 ;
    END
  END imonem
  PIN tmonem
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 54.3 7.1 54.5 7.3 ;
    END
  END tmonem
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER ME2 ;
        RECT 31.9 48.7 32.1 48.9 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 32.7 48.7 32.9 48.9 ;
    END
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 33.5 48.7 33.7 48.9 ;
    END
  END SO
  OBS
    LAYER ME1 SPACING 0.16 ;
      RECT 19.5 7.1 103.3 48.9 ;
    LAYER ME2 SPACING 0.2 ;
      RECT 34.06 7.66 103.3 48.9 ;
      RECT 54.86 7.1 103.3 48.9 ;
      RECT 19.5 7.66 31.54 48.9 ;
      RECT 24.06 7.1 39.54 48.34 ;
      RECT 53.66 7.1 53.94 48.9 ;
      RECT 52.46 7.1 52.74 48.9 ;
      RECT 51.26 7.1 51.54 48.9 ;
      RECT 47.26 7.1 47.54 48.9 ;
      RECT 43.26 7.1 43.54 48.9 ;
      RECT 22.46 7.1 23.14 48.9 ;
      RECT 19.5 7.1 20.74 48.9 ;
    LAYER ME3 SPACING 0.2 ;
      RECT 34 12.46 103.3 48.9 ;
      RECT 19.5 46.46 31.6 48.9 ;
      RECT 24 7.1 39.6 48.4 ;
      RECT 20.06 12.46 103.3 48.4 ;
      RECT 19.5 40.46 103.3 44.74 ;
      RECT 19.5 36.46 103.3 36.74 ;
      RECT 19.5 32.46 103.3 32.74 ;
      RECT 19.5 28.46 103.3 28.74 ;
      RECT 19.5 24.46 103.3 24.74 ;
      RECT 19.5 20.46 103.3 20.74 ;
      RECT 19.5 16.46 103.3 16.74 ;
      RECT 19.5 7.1 20.8 15.54 ;
      RECT 19.5 7.6 102.74 15.54 ;
      RECT 54.8 7.1 103.3 9.94 ;
      RECT 53.6 7.1 54 48.9 ;
      RECT 52.4 7.1 52.8 48.9 ;
      RECT 51.2 7.1 51.6 48.9 ;
      RECT 47.2 7.1 47.6 48.9 ;
      RECT 43.2 7.1 43.6 48.9 ;
      RECT 22.4 7.1 23.2 48.9 ;
    LAYER ME4 SPACING 0.2 ;
      RECT 19.5 46.4 103.3 48.9 ;
      RECT 20 12.4 103.3 48.9 ;
      RECT 19.5 40.4 103.3 44.8 ;
      RECT 19.5 36.4 103.3 36.8 ;
      RECT 19.5 32.4 103.3 32.8 ;
      RECT 19.5 28.4 103.3 28.8 ;
      RECT 19.5 24.4 103.3 24.8 ;
      RECT 19.5 20.4 103.3 20.8 ;
      RECT 19.5 16.4 103.3 16.8 ;
      RECT 19.5 7.1 102.8 15.6 ;
      RECT 19.5 7.1 103.3 10 ;
    LAYER ME5 SPACING 0.2 ;
      RECT 19.5 7.1 103.3 48.9 ;
    LAYER ME6 SPACING 0.2 ;
      RECT 19.5 7.1 103.3 48.9 ;
    LAYER ME7 SPACING 0.4 ;
      RECT 19.5 7.1 103.3 48.9 ;
    LAYER ME8 SPACING 1.5 ;
      RECT 19.5 7.1 103.3 48.9 ;
  END
END BATCHARGERctr

END LIBRARY